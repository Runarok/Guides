// 1. N-bit Decoder (2ⁿ to 2ⁿ outputs)
module decoder #(parameter N = 3) (
    input  wire [N-1:0] in,  // N-bit input signal
    output wire [(1<<N)-1:0] out  // 2ⁿ output signals
);
    // The decoder simply sets the output corresponding to the binary value of 'in'
    assign out = 1 << in;  // Left shift 1 by the value of 'in' to create the output
endmodule

//---

// 2. N-bit Multiplexer (2ⁿ inputs to 1 output)
module multiplexer #(parameter N = 3, WIDTH = 1) (
    input  wire [((1<<N)*WIDTH)-1:0] in,  // Concatenated inputs of size 2ⁿ * WIDTH
    input  wire [N-1:0] sel,  // N-bit select signal
    output wire [WIDTH-1:0] out  // 1-bit output (or WIDTH-bits if WIDTH > 1)
);
    // The multiplexer selects one of the inputs based on the value of 'sel'
    assign out = in[sel*WIDTH +: WIDTH];  // Use 'sel' to select the appropriate 'WIDTH' bits from 'in'
endmodule

//---

// 3. N-bit Binary to Gray Code Converter
module binary_to_gray #(parameter N = 4) (
    input  wire [N-1:0] bin,  // N-bit binary input
    output wire [N-1:0] gray  // N-bit Gray code output
);
    // The Gray code output is generated by XORing each bit of the input with its shifted version
    assign gray = bin ^ (bin >> 1);  // XOR the binary value with a right-shifted version of itself
endmodule

//---

// 4. N-bit Gray Code to Binary Converter
module gray_to_binary #(parameter N = 4) (
    input  wire [N-1:0] gray,  // N-bit Gray code input
    output reg  [N-1:0] bin  // N-bit binary output
);
    integer i;
    always @(*) begin
        // Start with the MSB (Most Significant Bit)
        bin[N-1] = gray[N-1];
        
        // Iterate through the rest of the bits to convert from Gray code to binary
        for (i = N-2; i >= 0; i = i - 1)
            bin[i] = bin[i+1] ^ gray[i];  // Perform XOR to reconstruct the binary number
    end
endmodule

//---

// 5. N-bit Binary Up-Down Counter
module up_down_counter #(parameter N = 4) (
    input  wire clk,  // Clock signal
    input  wire rst,  // Reset signal
    input  wire up_down,  // Control signal: 1 for counting up, 0 for counting down
    output reg  [N-1:0] count  // N-bit counter output
);
    always @(posedge clk or posedge rst) begin
        // Reset the counter to 0 on reset signal
        if (rst)
            count <= 0;
        // If counting up, increment the counter; if counting down, decrement it
        else if (up_down)
            count <= count + 1;
        else
            count <= count - 1;
    end
endmodule
