// Full Adder Module
// This module implements a 1-bit Full Adder, which takes in two input bits (A and B) 
// and a carry-in (Cin), producing a sum (S) and a carry-out (Cout).

module Full_Adder (
    input A,      // Input A (1-bit)
    input B,      // Input B (1-bit)
    input Cin,    // Carry-in (1-bit)
    output S,     // Sum output (1-bit)
    output Cout   // Carry-out output (1-bit)
);

// Sum is the result of the XOR operation between A, B, and Cin.
assign S = A ^ B ^ Cin;

// Carry-out is generated by checking if any two of the inputs are 1.
assign Cout = (A & B) | (B & Cin) | (Cin & A);

endmodule
