// megafunction wizard: %LPM_MULT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mult

// ============================================================
// File Name: MultiplyIP.v
// Megafunction Name(s): 
//             lpm_mult
//
// Simulation Library Files(s):
//             lpm
// ============================================================
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 24.1std.0 Build 1077 03/04/2025 SC Lite Edition
// ************************************************************

// Copyright (C) 2025  Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus Prime License Agreement,
// the Altera IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Altera and sold by Altera or its authorized distributors.  
// Please refer to the Altera Software License Subscription Agreements 
// on the Quartus Prime software download page.

// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on

module MultiplyIP (
    input   [7:0]  dataa,    // First input operand (8 bits)
    input   [7:0]  datab,    // Second input operand (8 bits)
    output  [15:0] result    // Output product (16 bits)
);

    // Internal wire for the result from the lpm_mult component
    wire [15:0] sub_wire0;
    wire [15:0] result = sub_wire0[15:0];

    // Instantiate the LPM_MULT component for multiplication
    lpm_mult lpm_mult_component (
        .dataa (dataa),           // Input operand A
        .datab (datab),           // Input operand B
        .result (sub_wire0),      // Result of multiplication
        .aclr (1'b0),             // Asynchronous clear (disabled)
        .clken (1'b1),            // Clock enable (enabled)
        .clock (1'b0),            // Clock (not used, set to 0)
        .sclr (1'b0),             // Synchronous clear (disabled)
        .sum (1'b0)               // Sum (not used, set to 0)
    );

    // Parameterize the LPM_MULT component with necessary settings
    defparam
        lpm_mult_component.lpm_hint               = "MAXIMIZE_SPEED=5", // Maximize speed optimization
        lpm_mult_component.lpm_representation     = "UNSIGNED",        // Unsigned multiplication
        lpm_mult_component.lpm_type               = "LPM_MULT",        // Use LPM_MULT megafunction
        lpm_mult_component.lpm_widtha             = 8,                 // Operand A width (8 bits)
        lpm_mult_component.lpm_widthb             = 8,                 // Operand B width (8 bits)
        lpm_mult_component.lpm_widthp             = 16;                // Product width (16 bits)

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
// Retrieval info: PRIVATE: ConstantB NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
// Retrieval info: PRIVATE: Latency NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SignedMult NUMERIC "0"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
// Retrieval info: PRIVATE: WidthA NUMERIC "8"
// Retrieval info: PRIVATE: WidthB NUMERIC "8"
// Retrieval info: PRIVATE: WidthP NUMERIC "16"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: PRIVATE: optimize NUMERIC "0"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=5"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
// Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "8"
// Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "8"
// Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "16"
// Retrieval info: USED_PORT: dataa 0 0 8 0 INPUT NODEFVAL "dataa[7..0]"
// Retrieval info: USED_PORT: datab 0 0 8 0 INPUT NODEFVAL "datab[7..0]"
// Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT NODEFVAL "result[15..0]"
// Retrieval info: CONNECT: @dataa 0 0 8 0 dataa 0 0 8 0
// Retrieval info: CONNECT: @datab 0 0 8 0 datab 0 0 8 0
// Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
// Retrieval info: GEN_FILE: TYPE_NORMAL MultiplyIP.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL MultiplyIP.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MultiplyIP.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MultiplyIP.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MultiplyIP_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL MultiplyIP_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
